/////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Mihai Olaru
// 
// Create Date: 02/18/2019 02:52:17 PM
// Design Name: Class with all the matrix computed
// Module Name: AlreadyComputed.sv
// Project Name: AES - Crypto
// Target Devices: 
// Tool Versions: 
// Description: aes_calculator
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
`include "ve_AES_types.sv"

`include "ve_AES_interface.sv"

`include "ve_AES_BaseUnit.sv"


`include "ve_AES_AlreadyComputed.sv"
`include "ve_AES_Core.sv"

//test_bench
`include "ve_AES_class_MixColumn.sv"

//`include "ve_AES_top_mix_column.sv"
`include "ve_AES_env.sv"