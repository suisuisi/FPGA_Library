/////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Mihai Olaru
// 
// Create Date: 02/18/2019 02:52:17 PM
// Design Name: Class with all the matrix computed
// Module Name: AlreadyComputed.sv
// Project Name: AES - Crypto
// Target Devices: 
// Tool Versions: 
// Description: aes_calculator
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`ifndef Cineva
`define Cineva
typedef bit [7 : 0]		word8;
typedef bit [31 : 0] word32;


`define 	MAXBC 8
`define 	MAXKC 8
`define  	MAXROUNDS 14
`define 	U_8 8
`endif