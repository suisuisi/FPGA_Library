/////////////////////////////
//   S-Box & Permutation   //
/////////////////////////////
module SP(S, P);
  input  [1:48] S;
  output [1:32] P;

  reg [1:4] x1, x2, x3, x4, x5, x6, x7, x8;

  assign P = {x4[4], x2[3], x5[4], x6[1], x8[1], x3[4], x7[4], x5[1],
              x1[1], x4[3], x6[3], x7[2], x2[1], x5[2], x8[3], x3[2],
              x1[2], x2[4], x6[4], x4[2], x8[4], x7[3], x1[3], x3[1],
              x5[3], x4[1], x8[2], x2[2], x6[2], x3[3], x1[4], x7[1]};

  always @(S[1:6]) begin
    case ({S[1], S[6], S[ 2: 5]})
       0: x1 =  9;   1: x1 =  7;   2: x1 = 15;   3: x1 =  2;
       4: x1 =  6;   5: x1 = 12;   6: x1 = 10;   7: x1 =  1;
       8: x1 =  3;   9: x1 =  0;  10: x1 =  4;  11: x1 = 14;
      12: x1 =  8;  13: x1 =  5;  14: x1 = 13;  15: x1 = 11;
      16: x1 =  3;  17: x1 =  0;  18: x1 =  5;  19: x1 = 11;
      20: x1 = 15;  21: x1 =  6;  22: x1 =  9;  23: x1 = 12;
      24: x1 =  8;  25: x1 = 13;  26: x1 =  2;  27: x1 =  4;
      28: x1 =  1;  29: x1 = 10;  30: x1 = 14;  31: x1 =  7;
      32: x1 =  6;  33: x1 = 10;  34: x1 =  0;  35: x1 =  7;
      36: x1 =  5;  37: x1 =  9;  38: x1 = 15;  39: x1 =  4;
      40: x1 = 12;  41: x1 =  3;  42: x1 = 11;  43: x1 =  8;
      44: x1 =  2;  45: x1 = 14;  46: x1 =  1;  47: x1 = 13;
      48: x1 = 15;  49: x1 =  6;  50: x1 = 10;  51: x1 =  0;
      52: x1 =  9;  53: x1 =  5;  54: x1 = 12;  55: x1 = 11;
      56: x1 =  2;  57: x1 =  8;  58: x1 =  1;  59: x1 = 13;
      60: x1 = 14;  61: x1 =  3;  62: x1 =  7;  63: x1 =  4;
    endcase
  end

  always @(S[7:12]) begin
    case ({S[7], S[12], S[ 8:11]})
       0: x2 =  8;   1: x2 =  4;   2: x2 =  2;   3: x2 =  9;
       4: x2 =  1;   5: x2 = 14;   6: x2 = 13;   7: x2 =  3;
       8: x2 =  5;   9: x2 = 11;  10: x2 = 15;  11: x2 = 12;
      12: x2 = 10;  13: x2 =  7;  14: x2 =  6;  15: x2 =  0;
      16: x2 = 15;  17: x2 =  1;  18: x2 =  5;  19: x2 = 10;
      20: x2 =  8;  21: x2 =  4;  22: x2 =  2;  23: x2 = 13;
      24: x2 =  9;  25: x2 =  7;  26: x2 =  6;  27: x2 =  0;
      28: x2 =  3;  29: x2 = 14;  30: x2 = 12;  31: x2 = 11;
      32: x2 = 14;  33: x2 =  3;  34: x2 =  4;  35: x2 = 15;
      36: x2 = 13;  37: x2 =  8;  38: x2 =  1;  39: x2 =  6;
      40: x2 =  0;  41: x2 =  5;  42: x2 =  9;  43: x2 =  2;
      44: x2 =  7;  45: x2 = 11;  46: x2 = 10;  47: x2 = 12;
      48: x2 =  0;  49: x2 = 13;  50: x2 = 14;  51: x2 =  4;
      52: x2 = 11;  53: x2 =  1;  54: x2 =  7;  55: x2 = 10;
      56: x2 =  6;  57: x2 =  8;  58: x2 =  3;  59: x2 = 15;
      60: x2 = 12;  61: x2 =  2;  62: x2 =  9;  63: x2 =  5;
    endcase
  end

  always @(S[13:18]) begin
    case ({S[13], S[18], S[14:17]})
       0: x3 = 14;   1: x3 =  3;   2: x3 =  4;   3: x3 = 15;
       4: x3 =  2;   5: x3 = 12;   6: x3 = 11;   7: x3 =  5;
       8: x3 = 13;   9: x3 =  0;  10: x3 =  1;  11: x3 = 10;
      12: x3 =  8;  13: x3 =  7;  14: x3 =  6;  15: x3 =  9;
      16: x3 =  2;  17: x3 = 12;  18: x3 = 11;  19: x3 =  1;
      20: x3 = 14;  21: x3 =  7;  22: x3 =  5;  23: x3 = 10;
      24: x3 =  4;  25: x3 =  9;  26: x3 = 13;  27: x3 =  6;
      28: x3 =  3;  29: x3 =  0;  30: x3 =  8;  31: x3 = 15;
      32: x3 =  5;  33: x3 = 14;  34: x3 =  2;  35: x3 =  8;
      36: x3 = 15;  37: x3 =  1;  38: x3 = 12;  39: x3 = 11;
      40: x3 =  0;  41: x3 =  9;  42: x3 = 13;  43: x3 =  7;
      44: x3 =  6;  45: x3 = 10;  46: x3 =  3;  47: x3 =  4;
      48: x3 = 12;  49: x3 =  7;  50: x3 =  1;  51: x3 = 13;
      52: x3 =  2;  53: x3 =  8;  54: x3 = 11;  55: x3 =  4;
      56: x3 =  9;  57: x3 = 14;  58: x3 = 10;  59: x3 =  0;
      60: x3 = 15;  61: x3 =  5;  62: x3 =  6;  63: x3 =  3;
    endcase
  end

  always @(S[19:24]) begin
    case ({S[19], S[24], S[20:23]})
       0: x4 = 13;   1: x4 =  3;   2: x4 =  6;   3: x4 =  5;
       4: x4 =  8;   5: x4 = 15;   6: x4 = 11;   7: x4 =  0;
       8: x4 =  4;   9: x4 = 10;  10: x4 =  9;  11: x4 = 12;
      12: x4 =  2;  13: x4 =  1;  14: x4 = 14;  15: x4 =  7;
      16: x4 =  4;  17: x4 =  9;  18: x4 =  3;  19: x4 =  0;
      20: x4 = 14;  21: x4 =  5;  22: x4 = 13;  23: x4 = 10;
      24: x4 =  2;  25: x4 = 15;  26: x4 = 12;  27: x4 =  6;
      28: x4 = 11;  29: x4 =  8;  30: x4 =  7;  31: x4 =  1;
      32: x4 = 10;  33: x4 =  4;  34: x4 =  5;  35: x4 =  8;
      36: x4 = 15;  37: x4 =  3;  38: x4 =  6;  39: x4 = 13;
      40: x4 =  7;  41: x4 =  1;  42: x4 = 14;  43: x4 =  2;
      44: x4 =  9;  45: x4 = 12;  46: x4 =  0;  47: x4 = 11;
      48: x4 = 15;  49: x4 =  2;  50: x4 =  0;  51: x4 = 14;
      52: x4 =  5;  53: x4 =  9;  54: x4 =  3;  55: x4 =  4;
      56: x4 =  1;  57: x4 =  8;  58: x4 =  7;  59: x4 = 11;
      60: x4 = 12;  61: x4 =  6;  62: x4 = 10;  63: x4 = 13;
    endcase
  end

  always @(S[25:30]) begin
    case ({S[25], S[30], S[26:29]})
       0: x5 =  8;   1: x5 =  6;   2: x5 =  7;   3: x5 =  1;
       4: x5 =  4;   5: x5 = 13;   6: x5 =  2;   7: x5 = 11;
       8: x5 =  3;   9: x5 = 12;  10: x5 =  0;  11: x5 = 15;
      12: x5 =  9;  13: x5 = 10;  14: x5 = 14;  15: x5 =  5;
      16: x5 =  4;  17: x5 =  1;  18: x5 =  2;  19: x5 = 12;
      20: x5 = 13;  21: x5 = 11;  22: x5 = 14;  23: x5 =  7;
      24: x5 =  8;  25: x5 = 15;  26: x5 =  5;  27: x5 = 10;
      28: x5 =  6;  29: x5 =  0;  30: x5 =  3;  31: x5 =  9;
      32: x5 =  1;  33: x5 = 11;  34: x5 = 10;  35: x5 =  4;
      36: x5 =  7;  37: x5 =  2;  38: x5 = 13;  39: x5 =  8;
      40: x5 =  6;  41: x5 =  5;  42: x5 = 15;  43: x5 =  3;
      44: x5 = 12;  45: x5 =  9;  46: x5 =  0;  47: x5 = 14;
      48: x5 = 15;  49: x5 =  2;  50: x5 = 12;  51: x5 = 11;
      52: x5 = 10;  53: x5 =  7;  54: x5 =  1;  55: x5 = 13;
      56: x5 =  5;  57: x5 =  8;  58: x5 =  9;  59: x5 =  4;
      60: x5 =  0;  61: x5 = 14;  62: x5 =  6;  63: x5 =  3;
    endcase
  end

  always @(S[31:36]) begin
    case ({S[31], S[36], S[32:35]})
       0: x6 = 15;   1: x6 =  4;   2: x6 = 12;   3: x6 =  7;
       4: x6 =  5;   5: x6 =  2;   6: x6 = 10;   7: x6 =  9;
       8: x6 =  8;   9: x6 =  3;  10: x6 =  1;  11: x6 = 13;
      12: x6 = 11;  13: x6 = 14;  14: x6 =  6;  15: x6 =  0;
      16: x6 =  3;  17: x6 = 10;  18: x6 = 15;  19: x6 =  1;
      20: x6 =  9;  21: x6 =  4;  22: x6 =  0;  23: x6 =  7;
      24: x6 =  6;  25: x6 = 13;  26: x6 = 12;  27: x6 =  2;
      28: x6 =  5;  29: x6 =  8;  30: x6 = 11;  31: x6 = 14;
      32: x6 =  4;  33: x6 =  2;  34: x6 =  9;  35: x6 = 12;
      36: x6 = 10;  37: x6 = 15;  38: x6 =  3;  39: x6 =  5;
      40: x6 =  1;  41: x6 = 13;  42: x6 = 14;  43: x6 = 11;
      44: x6 =  7;  45: x6 =  0;  46: x6 =  8;  47: x6 =  6;
      48: x6 =  9;  49: x6 =  5;  50: x6 =  2;  51: x6 = 15;
      52: x6 =  4;  53: x6 =  3;  54: x6 = 14;  55: x6 =  0;
      56: x6 = 12;  57: x6 =  6;  58: x6 =  7;  59: x6 =  8;
      60: x6 = 10;  61: x6 = 13;  62: x6 =  1;  63: x6 = 11;
    endcase
  end

  always @(S[37:42]) begin
    case ({S[37], S[42], S[38:41]})
       0: x7 =  3;   1: x7 = 12;   2: x7 = 14;   3: x7 =  2;
       4: x7 =  0;   5: x7 = 15;   6: x7 =  9;   7: x7 =  5;
       8: x7 = 10;   9: x7 =  7;  10: x7 =  1;  11: x7 =  4;
      12: x7 = 13;  13: x7 =  8;  14: x7 =  6;  15: x7 = 11;
      16: x7 =  9;  17: x7 =  2;  18: x7 =  0;  19: x7 =  5;
      20: x7 =  6;  21: x7 =  8;  22: x7 = 10;  23: x7 = 15;
      24: x7 =  7;  25: x7 = 14;  26: x7 = 12;  27: x7 =  3;
      28: x7 = 11;  29: x7 = 13;  30: x7 =  1;  31: x7 =  4;
      32: x7 =  8;  33: x7 =  6;  34: x7 =  2;  35: x7 = 15;
      36: x7 =  5;  37: x7 = 12;  38: x7 = 14;  39: x7 =  3;
      40: x7 =  1;  41: x7 = 10;  42: x7 =  4;  43: x7 =  9;
      44: x7 = 11;  45: x7 =  7;  46: x7 = 13;  47: x7 =  0;
      48: x7 =  6;  49: x7 =  1;  50: x7 =  5;  51: x7 = 10;
      52: x7 =  9;  53: x7 =  7;  54: x7 =  3;  55: x7 = 12;
      56: x7 =  8;  57: x7 = 13;  58: x7 = 15;  59: x7 =  0;
      60: x7 =  2;  61: x7 = 14;  62: x7 =  4;  63: x7 = 11;
    endcase
  end

  always @(S[43:48]) begin
    case ({S[43], S[48], S[44:47]})
       0: x8 = 11;   1: x8 =  0;   2: x8 =  7;   3: x8 =  9;
       4: x8 =  2;   5: x8 = 15;   6: x8 = 12;   7: x8 =  5;
       8: x8 = 13;   9: x8 = 14;  10: x8 = 10;  11: x8 =  3;
      12: x8 =  1;  13: x8 =  4;  14: x8 =  6;  15: x8 =  8;
      16: x8 = 14;  17: x8 =  5;  18: x8 =  9;  19: x8 = 12;
      20: x8 =  7;  21: x8 = 10;  22: x8 =  0;  23: x8 =  3;
      24: x8 =  8;  25: x8 =  2;  26: x8 =  6;  27: x8 = 15;
      28: x8 = 13;  29: x8 =  1;  30: x8 = 11;  31: x8 =  4;
      32: x8 =  2;  33: x8 = 15;  34: x8 = 12;  35: x8 = 10;
      36: x8 =  9;  37: x8 =  0;  38: x8 =  5;  39: x8 =  6;
      40: x8 =  4;  41: x8 =  1;  42: x8 =  3;  43: x8 = 13;
      44: x8 = 14;  45: x8 =  7;  46: x8 =  8;  47: x8 = 11;
      48: x8 =  1;  49: x8 = 12;  50: x8 = 10;  51: x8 =  6;
      52: x8 =  4;  53: x8 =  3;  54: x8 = 15;  55: x8 =  9;
      56: x8 = 11;  57: x8 =  7;  58: x8 =  5;  59: x8 =  0;
      60: x8 =  8;  61: x8 = 13;  62: x8 =  2;  63: x8 = 14;
    endcase
  end
endmodule


/////////////////////////////
//         DES core        //
/////////////////////////////
module DES(Din, Key, Dout, Drdy, Krdy, ENC, RSTn, EN, CLK, BSY, Dvld);
  input  [1:64] Din;  // Data input
  input  [1:64] Key;  // Key input
  output [1:64] Dout; // Data output
  input  Drdy;        // Data input ready
  input  Krdy;        // Key input ready
  input  ENC;         // 1 encryption, 0 decryption
  input  RSTn;        // Reset (Low active)
  input  EN;          // DES circuit enable
  input  CLK;         // System clock
  output BSY;         // Busy signal
  output Dvld;        // Data output valid

  reg  [1:64] Drg;    // Data register
  reg  [1:56] Krg;    // Key Register
  reg  [1:16] Rrg;    // Round Register
  reg  BSYrg;         // 0 WAIT, 1 ROUND (busy)
  reg  Dvldrg;

  wire [1:64] Mask;
  wire [1:32] MaskLR;
  wire [1:64] DiX, DoX;
  wire [1:64] IP;
  wire [1:56] PC1, PC2, Knext;
  wire [1:48] Kadd, Sin;
  wire [1:32] Pout;

  assign Mask   = 64'h0123456789abcdef;
  assign MaskLR = Mask[1:32] ^ Mask[33:64];
  assign DiX   = IP ^ Mask;
  assign DoX   = Drg ^ Mask;
 
  assign IP   = {Din[58], Din[50], Din[42], Din[34], Din[26], Din[18], Din[10], Din[2],
                 Din[60], Din[52], Din[44], Din[36], Din[28], Din[20], Din[12], Din[4],
                 Din[62], Din[54], Din[46], Din[38], Din[30], Din[22], Din[14], Din[6],
                 Din[64], Din[56], Din[48], Din[40], Din[32], Din[24], Din[16], Din[8],
                 Din[57], Din[49], Din[41], Din[33], Din[25], Din[17], Din[ 9], Din[1],
                 Din[59], Din[51], Din[43], Din[35], Din[27], Din[19], Din[11], Din[3],
                 Din[61], Din[53], Din[45], Din[37], Din[29], Din[21], Din[13], Din[5],
                 Din[63], Din[55], Din[47], Din[39], Din[31], Din[23], Din[15], Din[7]};

  assign Dout = {DoX[8], DoX[40], DoX[16], DoX[48], DoX[24], DoX[56], DoX[32], DoX[64],
                 DoX[7], DoX[39], DoX[15], DoX[47], DoX[23], DoX[55], DoX[31], DoX[63],
                 DoX[6], DoX[38], DoX[14], DoX[46], DoX[22], DoX[54], DoX[30], DoX[62],
                 DoX[5], DoX[37], DoX[13], DoX[45], DoX[21], DoX[53], DoX[29], DoX[61],
                 DoX[4], DoX[36], DoX[12], DoX[44], DoX[20], DoX[52], DoX[28], DoX[60],
                 DoX[3], DoX[35], DoX[11], DoX[43], DoX[19], DoX[51], DoX[27], DoX[59],
                 DoX[2], DoX[34], DoX[10], DoX[42], DoX[18], DoX[50], DoX[26], DoX[58],
                 DoX[1], DoX[33], DoX[ 9], DoX[41], DoX[17], DoX[49], DoX[25], DoX[57]};

  assign PC1  = {Key[57], Key[49], Key[41], Key[33], Key[25], Key[17], Key[ 9],
                 Key[ 1], Key[58], Key[50], Key[42], Key[34], Key[26], Key[18],
                 Key[10], Key[ 2], Key[59], Key[51], Key[43], Key[35], Key[27],
                 Key[19], Key[11], Key[ 3], Key[60], Key[52], Key[44], Key[36],
                 Key[63], Key[55], Key[47], Key[39], Key[31], Key[23], Key[15],
                 Key[ 7], Key[62], Key[54], Key[46], Key[38], Key[30], Key[22],
                 Key[14], Key[ 6], Key[61], Key[53], Key[45], Key[37], Key[29],
                 Key[21], Key[13], Key[ 5], Key[28], Key[20], Key[12], Key[ 4]};

  assign Knext = (ENC == 1)? 
                 (((Rrg[1] | Rrg[2] | Rrg[9] | Rrg[16]) == 1)?
                   {Krg[2:28], Krg[1], Krg[30:56], Krg[29]}:
                   {Krg[3:28], Krg[1:2], Krg[31:56], Krg[29:30]}):
                 (((Rrg[1] | Rrg[8] | Rrg[15] | Rrg[16]) == 1)?
                   {Krg[28], Krg[1:27], Krg[56], Krg[29:55]}:
                   {Krg[27:28], Krg[1:26], Krg[55:56], Krg[29:54]});

  assign PC2 = (ENC ==1)? Knext: Krg;
  assign Kadd = {PC2[14], PC2[17], PC2[11], PC2[24], PC2[ 1], PC2[ 5],
                 PC2[ 3], PC2[28], PC2[15], PC2[ 6], PC2[21], PC2[10],
                 PC2[23], PC2[19], PC2[12], PC2[ 4], PC2[26], PC2[ 8],
                 PC2[16], PC2[ 7], PC2[27], PC2[20], PC2[13], PC2[ 2],
                 PC2[41], PC2[52], PC2[31], PC2[37], PC2[47], PC2[55],
                 PC2[30], PC2[40], PC2[51], PC2[45], PC2[33], PC2[48],
                 PC2[44], PC2[49], PC2[39], PC2[56], PC2[34], PC2[53],
                 PC2[46], PC2[42], PC2[50], PC2[36], PC2[29], PC2[32]};

  assign Sin = {Drg[64], Drg[33:37], Drg[36:41], Drg[40:45], Drg[44:49],
                Drg[48:53], Drg[52:57], Drg[56:61], Drg[60:64], Drg[33]} ^ Kadd;
  SP SP (Sin, Pout);

  assign BSY = BSYrg;
  assign Dvld = Dvldrg;

  always @(posedge CLK) begin
    if (RSTn == 0) begin
       Rrg    <= 16'b1000000000000000;
       BSYrg  <= 0;
       Dvldrg <= 0;
    end
    else if (EN == 1) begin
      if (BSYrg == 0) begin  // Idol
        if (Krdy == 1)
          Krg <= PC1;
        if (Drdy == 1) begin
          BSYrg  <= 1;
          Drg    <= DiX;
          Dvldrg <= 0;
        end
      end
      else begin  // Round
        Drg <= {Drg[33:64] ^ MaskLR, Drg[1:32] ^ Pout};
        Krg <= Knext;
        Rrg <= {Rrg[16], Rrg[1:15]};
        if (Rrg[16] == 1) begin
          BSYrg  <= 0;
          Dvldrg <= 1;
        end
      end
    end
  end
endmodule
